* ADG849 SPICE Macro-model
* Generic Desc: 0.35 CMOS 1.65 V to 3.6 V Single SPDT Switch/2:1 MUX
* Developed by: MPorley / ADGT
* Revision History: 1.0 (8/2018)
* Copyright 2018 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model
* indicates your acceptance of the terms and provisions in the License Statement.
*
* Begin Notes:
* The model will work on Vdd/Vss from 1.65V to 3.6V single supply.
* The model provides parametric specifications at +3.6V only and is not variable with Vdd. Please see datasheet page 3.
*
* Not Modeled:
*
* Parameters modeled include:
*	On Resistance
*	Ton and Toff
*	Break-Before-Make
*	Off Isolation
*	Crosstalk
*	Supply Currents: Iss/Idd
*	Bandwidth
*	Charge Injection
* Connections
*      1  = IN1
*      2  = VDD
*      3  = GND
*      4  = S1
*      5  = D1
*      6  = S2
*
.SUBCKT ADG849 1 2 3 4 5 6

.MODEL VON VSWITCH(Von=5 Voff=0.8 Ron=0.001 Roff=1000000000000)
.MODEL VEN VSWITCH(Von=5 Voff=0.8 Ron=12000 Roff=21000)
.MODEL VNE VSWITCH(Von=5 Voff=0.8 Ron=14000 Roff=11000)
.MODEL VRESET VSWITCH(Von=5 Voff=0.8 Ron=2700000 Roff=1000)
.MODEL DCLAMP D(IS=1E-15 IBV=1E-13)


* CROSSTALK
C12X 4 6 3.8E-012

* IDD/ISS
I1 2 3 0.003E-006

* Configuration: SPST 2:2


** SWITCH 1 **
*
* ESD PROTECTION DIODES
D11 3 5 DCLAMP
D12 5 2 DCLAMP
D13 3 4 DCLAMP
D14 4 2 DCLAMP
*
* OFF ISOLATION
C11 4 5 3.8E-012
*
* CHARGE INJECTION
C12 5 140 2.5E-011
C13 4 140 2.5E-011
*
* CD/CS OFF AND BANDWIDTH
C14 4 3 90E-012
C15 5 3 75e-012
*
* ON RESISTANCE
Ech155 1555 3 VALUE = { IF ((ABS(V(4)))>(ABS(V(184))),V(4),V(5)) }
R155 1555 3 1G
R11 137 5 0.001
S111 136 141 1141 3 VON
Ech111 1141 3 VALUE = { IF (V(1555)<1,5,0) }
Ech11 141 3 VALUE = { IF (V(1555)<1,0.01*(V(1555)-1)+0.34,0) }
S112 136 146 1146 3 VON
Ech112 1146 3 VALUE = { IF ((V(1555)>=1) & (V(1555)<=2.7),5,0) }
Ech12 146 3 VALUE = { IF ((V(1555)>=1) & (V(1555)<=2.7),((0.34-0.28)/((1-1.9358674372686)*(1-1.9358674372686)))*(V(1555)-1.9358674372686)*(V(1555)-1.9358674372686) + 0.28,0) }
S113 136 144 1144 3 VON
Ech113 1144 3 VALUE = { IF (V(1555)>2.7,5,0) }
Ech13 144 3 VALUE = { IF (V(1555)>2.7,-1.11111111111111E-02*(V(1555)-2.7)+0.32,0) }
RIN1	136 3	1G
EOUT1 137 181	POLY(2) (136,3) (180,3) 0 0 0 0 0.999/1000
FCOPY1	3 180 VSENSE1 1
RSENSOR1 180 3	1K
VSENSE1 181 184	0
*
* TON/ TOFF/ BBM
S11 182 184 140 3 VON
S12 143 138 143 3 VEN
Ech14 143 3 VALUE = { IF(V(1)>=2.0, 5 , 0.8 ) }
eV1 140 3 138 3 1
C16 138 3 1e-012
*
* VOLTAGE SUPPLY REQUIREMENT
S13 4 182 185 3 VON
S15 139 185 139 3 VON
Ech16 139 3 VALUE = { IF((V(3)>=-0.5 & (V(2)<=3.6 & V(2)>=1.65)), 5 , 0.01 ) }


** SWITCH 2 **
*
* ESD PROTECTION DIODES
D21 3 7 DCLAMP
D22 7 2 DCLAMP
D23 3 6 DCLAMP
D24 6 2 DCLAMP
*
* OFF ISOLATION
C21 6 7 3.8E-012
*
* CHARGE INJECTION
C22 7 240 2.5E-011
C23 6 240 2.5E-011
*
* CD/CS OFF AND BANDWIDTH
C24 6 3 90E-012
C25 7 3 75e-012
*
* ON RESISTANCE
Ech255 2555 3 VALUE = { IF ((ABS(V(6)))>(ABS(V(284))),V(6),V(7)) }
R255 2555 3 1G
R21 237 5 0.001
S221 236 241 2241 3 VON
Ech221 2241 3 VALUE = { IF (V(2555)<1,5,0) }
Ech21 241 3 VALUE = { IF (V(2555)<1,0.01*(V(2555)-1)+0.34,0) }
S222 236 246 2246 3 VON
Ech222 2246 3 VALUE = { IF ((V(2555)>=1) & (V(2555)<=2.7),5,0) }
Ech22 246 3 VALUE = { IF ((V(2555)>=1) & (V(2555)<=2.7),((0.34-0.28)/((1-1.9358674372686)*(1-1.9358674372686)))*(V(2555)-1.9358674372686)*(V(2555)-1.9358674372686) + 0.28,0) }
S223 236 244 2244 3 VON
Ech223 2244 3 VALUE = { IF (V(2555)>2.7,5,0) }
Ech23 244 3 VALUE = { IF (V(2555)>2.7,-1.11111111111111E-02*(V(2555)-2.7)+0.32,0) }
RIN2	236 3	1G
EOUT2 237 281	POLY(2) (236,3) (280,3) 0 0 0 0 0.999/1000
FCOPY2	3 280 VSENSE2 1
RSENSOR2 280 3	1K
VSENSE2 281 284	0
*
* TON/ TOFF/ BBM
S21 282 284 240 3 VON
S22 243 238 243 3 VNE
Ech24 243 3 VALUE = { IF(V(1)<2.0, 5 , 0.8 ) }
eV2 240 3 238 3 1
C26 238 3 1e-012
*
* VOLTAGE SUPPLY REQUIREMENT
S23 6 282 285 3 VON
S25 239 285 239 3 VON
Ech26 239 3 VALUE = { IF((V(3)>=-0.5 & (V(2)<=3.6 & V(2)>=1.65)), 5 , 0.01 ) }

.ENDS ADG849
